`ifndef __INTERFACE_SV__
`define __INTERFACE_SV__

interface my_interface(output [31:0] foo);
endinterface

`endif
