interface ifc;
    logic val;
    byte  x;
endinterface
