`include "uvm_unit.svh"
import uvm_unit_pkg::*;

// Nothing here
