`include "fixtures_and_assertions_test.sv"
`include "second_file_test.sv"
